
`timescale 1ns / 1ps
`include "defines.sv"

module DataPath (
    //global signals
    input logic clk,
    input logic reset,

    // instruction memory side port
    input  logic [31:0] instrCode,
    output logic [31:0] instrMemAddr,

    //control unit side port
    input logic       PCEn,
    input logic       regFileWe,
    input logic [3:0] aluControl,
    input logic       aluSrcMuxSel,
    input logic [2:0] RFWDSrcMuxSel,
    input logic       branch,
    input logic       jal,
    input logic       jalr,

    //data memory side port
    output logic [31:0] busAddr,
    output logic [31:0] busWData,
    input  logic [31:0] busRData
);

    logic [31:0] aluResult, ExeReg_aluResult, RFData1, RFData2;
    logic [31:0] DecReg_RFData1, DecReg_RFData2, ExeReg_RFData2;
    logic [31:0] PCSrcData, PCOutData, PC_Imm_AdderSrcMuxOut;
    logic [31:0] aluSrcMuxOut, immExt, DecReg_immExt, RFWDSrcMuxOut;
    logic [31:0]
        PC_4_AdderResult, PC_Imm_AdderResult, PCSrcMuxOut, ExeReg_PCSrcMuxOut;
    logic [31:0] MemAccReg_busRData, LoadExtData, ConcatData;
    logic PCSrcMuxSel;
    logic btaken;

    assign instrMemAddr = PCOutData;
    assign busAddr = ExeReg_aluResult;
    assign busWData = ConcatData;

    RegisterFile U_RegFile (
        .clk(clk),
	.reset(reset),
        .we (regFileWe),
        .RA1(instrCode[19:15]),
        .RA2(instrCode[24:20]),
        .WA (instrCode[11:7]),
        .WD (RFWDSrcMuxOut),
        .RD1(RFData1),
        .RD2(RFData2)
    );

    data_extension_load LOAD_EXT (  //mem access operation
        .instrCode(instrCode),
        .busRData(busRData),
        .addr(ExeReg_aluResult),
        .ext_data(LoadExtData)
    );

    store_bit_concat STORE_CONCAT (  //mem access operation
        .instrCode(instrCode),
        .RFData2(ExeReg_RFData2),
        .busRData(busRData),
        .addr(ExeReg_aluResult),
        .concat_data(ConcatData)
    );

    register U_DecReg_RFRD1 (
        .clk(clk),
        .reset(reset),
        .d(RFData1),
        .q(DecReg_RFData1)
    );

    register U_DecReg_RFRD2 (
        .clk(clk),
        .reset(reset),
        .d(RFData2),
        .q(DecReg_RFData2)
    );

    register U_ExeReg_RFRD2 (
        .clk(clk),
        .reset(reset),
        .d(DecReg_RFData2),
        .q(ExeReg_RFData2)
    );

    register U_DecReg_ImmExtend (
        .clk(clk),
        .reset(reset),
        .d(immExt),
        .q(DecReg_immExt)
    );

    mux_2x1 U_AluSrcMux (
        .sel(aluSrcMuxSel),
        .x0 (DecReg_RFData2),
        .x1 (DecReg_immExt),
        .y  (aluSrcMuxOut)
    );

    register U_MemAccReg_ReadData (
        .clk(clk),
        .reset(reset),
        .d(LoadExtData),
        .q(MemAccReg_busRData)
    );

    mux_5x1 U_RFWDSrcMux (
        .sel(RFWDSrcMuxSel),
        .x0 (aluResult),
        .x1 (MemAccReg_busRData),
        .x2 (DecReg_immExt),
        .x3 (PC_Imm_AdderResult),
        .x4 (PC_4_AdderResult),
        .y  (RFWDSrcMuxOut)
    );

    alu U_ALU (
        .aluControl(aluControl),
        .a         (DecReg_RFData1),
        .b         (aluSrcMuxOut),
        .result    (aluResult),
        .btaken    (btaken)
    );

    register U_ExeReg_ALU (
        .clk(clk),
        .reset(reset),
        .d(aluResult),
        .q(ExeReg_aluResult)
    );

    immExtend U_ImmExtend (
        .instrCode(instrCode),
        .immExt   (immExt)
    );

    mux_2x1 U_PC_Imm_AdderSrcMux (
        .sel(jalr),
        .x0 (PCOutData),
        .x1 (DecReg_RFData1),
        .y  (PC_Imm_AdderSrcMuxOut)
    );

    adder U_PC_Imm_Adder (
        .a(DecReg_immExt),
        .b(PC_Imm_AdderSrcMuxOut),
        .y(PC_Imm_AdderResult)
    );

    adder U_PC_4_Adder (
        .a(32'd4),
        .b(PCOutData),
        .y(PC_4_AdderResult)
    );

    assign PCSrcMuxSel = jal | (btaken & branch);

    mux_2x1 U_PCSrcMux (
        .sel(PCSrcMuxSel),
        .x0 (PC_4_AdderResult),
        .x1 (PC_Imm_AdderResult),
        .y  (PCSrcMuxOut)
    );

    register U_ExeReg_PCSrcMux (
        .clk(clk),
        .reset(reset),
        .d(PCSrcMuxOut),
        .q(ExeReg_PCSrcMuxOut)
    );

    registerEn U_PC (
        .clk  (clk),
        .reset(reset),
        .en   (PCEn),
        .d    (ExeReg_PCSrcMuxOut),
        .q    (PCOutData)
    );

endmodule

module alu (
    input  logic [ 3:0] aluControl,
    input  logic [31:0] a,
    input  logic [31:0] b,
    output logic [31:0] result,
    output logic        btaken
);

    always_comb begin
        result = 32'bx;
        case (aluControl)
            `ADD:  result = a + b;
            `SUB:  result = a - b;
            `SLL:  result = a << b;
            `SRL:  result = a >> b;
            `SRA:  result = $signed(a) >>> b;
            `SLT:  result = ($signed(a) < $signed(b)) ? 1 : 0;
            `SLTU: result = (a < b) ? 1 : 0;
            `XOR:  result = a ^ b;
            `OR:   result = a | b;
            `AND:  result = a & b;
        endcase
    end

    always_comb begin : branch
        btaken = 1'b0;
        case (aluControl[2:0])
            `BEQ:  btaken = (a == b);
            `BNE:  btaken = (a != b);
            `BLT:  btaken = ($signed(a) < $signed(b));
            `BGE:  btaken = ($signed(a) >= $signed(b));
            `BLTU: btaken = (a < b);
            `BGEU: btaken = (a >= b);
        endcase
    end
endmodule


module RegisterFile (
    input  logic        clk,
    input  logic        reset,    // reset 추가
    input  logic        we,
    input  logic [ 4:0] RA1,
    input  logic [ 4:0] RA2,
    input  logic [ 4:0] WA,
    input  logic [31:0] WD,
    output logic [31:0] RD1,
    output logic [31:0] RD2
);
    logic [31:0] mem[0:31];



    // 초기값 할당: x0~x31
    always_ff @(posedge clk, posedge reset) begin
        if (reset) begin
            for (int i = 0; i < 32; i=i+1) begin
                if (i == 0)
                    mem[i] <= 32'd0;        // x0 항상 0
                else
                    mem[i] <= 9 + i;  // x1=10, x2=11, ..., x31=40
            end
        end else if (we && WA != 0) begin
            mem[WA] <= WD;
        end
    end

    assign RD1 = (RA1 != 0) ? mem[RA1] : 32'd0;
    assign RD2 = (RA2 != 0) ? mem[RA2] : 32'd0;

endmodule


module registerEn (
    input  logic        clk,
    input  logic        reset,
    input  logic        en,
    input  logic [31:0] d,
    output logic [31:0] q
);
    always_ff @(posedge clk, posedge reset) begin
        if (reset) begin
            q <= 0;
        end else begin
            if (en) q <= d;
        end
    end
endmodule

module register (
    input  logic        clk,
    input  logic        reset,
    input  logic [31:0] d,
    output logic [31:0] q
);
    always_ff @(posedge clk, posedge reset) begin
        if (reset) begin
            q <= 0;
        end else begin
            q <= d;
        end
    end
endmodule

module adder (
    input  logic [31:0] a,
    input  logic [31:0] b,
    output logic [31:0] y
);
    assign y = a + b;
endmodule

module mux_2x1 (
    input  logic        sel,
    input  logic [31:0] x0,
    input  logic [31:0] x1,
    output logic [31:0] y
);
    always_comb begin
        y = 32'bx;
        case (sel)
            1'b0: y = x0;
            1'b1: y = x1;
        endcase
    end
endmodule

module mux_5x1 (
    input  logic [ 2:0] sel,
    input  logic [31:0] x0,
    input  logic [31:0] x1,
    input  logic [31:0] x2,
    input  logic [31:0] x3,
    input  logic [31:0] x4,
    output logic [31:0] y
);
    always_comb begin
        y = 32'bx;
        case (sel)
            3'b000: y = x0;
            3'b001: y = x1;
            3'b010: y = x2;
            3'b011: y = x3;
            3'b100: y = x4;
        endcase
    end
endmodule

module immExtend (
    input  logic [31:0] instrCode,
    output logic [31:0] immExt
);
    wire [6:0] opcode = instrCode[6:0];
    wire [2:0] func3 = instrCode[14:12];

    always_comb begin
        immExt = 32'bx;
        case (opcode)
            `OP_TYPE_R: immExt = 32'bx;  // R-Type
            `OP_TYPE_L: immExt = {{20{instrCode[31]}}, instrCode[31:20]};
            `OP_TYPE_S:
            immExt = {
                {20{instrCode[31]}}, instrCode[31:25], instrCode[11:7]
            };  // S-Type
            `OP_TYPE_I: begin
                case (func3)
                    3'b001:  immExt = {27'b0, instrCode[24:20]};  // SLLI
                    3'b101:  immExt = {27'b0, instrCode[24:20]};  // SRLI, SRAI
                    3'b011:  immExt = {20'b0, instrCode[31:20]};  // SLTIU
                    default: immExt = {{20{instrCode[31]}}, instrCode[31:20]};
                endcase
            end
            `OP_TYPE_B:
            immExt = {
                {20{instrCode[31]}},
                instrCode[7],
                instrCode[30:25],
                instrCode[11:8],
                1'b0
            };
            `OP_TYPE_LU: immExt = {instrCode[31:12], 12'b0};
            `OP_TYPE_AU: immExt = {instrCode[31:12], 12'b0};
            `OP_TYPE_J:
            immExt = {
                {12{instrCode[31]}},
                instrCode[19:12],
                instrCode[20],
                instrCode[30:21],
                1'b0
            };
            `OP_TYPE_JL: immExt = {{20{instrCode[31]}}, instrCode[31:20]};
        endcase
    end
endmodule



module data_extension_load (
    input  logic [31:0] instrCode,
    input  logic [31:0] busRData,
    input  logic [31:0] addr,
    output logic [31:0] ext_data
);

    wire [6:0] opcode = instrCode[6:0];
    wire [2:0] func3 = instrCode[14:12];
    wire [1:0] byte_remain = addr[1:0];
    wire half_remain = addr[1];




    always_comb begin
        ext_data = 32'bx;
        case (opcode)
            `OP_TYPE_L: begin
                case (func3)
                    3'b000: begin
                        case (byte_remain)
                            2'b00:
                            ext_data = {{24{busRData[7]}}, busRData[7:0]};
                            2'b01:
                            ext_data = {{24{busRData[15]}}, busRData[15:8]};
                            2'b10:
                            ext_data = {{24{busRData[23]}}, busRData[23:16]};
                            2'b11:
                            ext_data = {{24{busRData[31]}}, busRData[31:24]};
                        endcase
                    end
                    3'b001: begin
                        case (half_remain)
                            0: ext_data = {{16{busRData[15]}}, busRData[15:0]};
                            1: ext_data = {{16{busRData[31]}}, busRData[31:16]};
                        endcase
                    end
                    3'b010: begin
                        ext_data = busRData;
                    end
                    3'b100: begin
                        case (byte_remain)
                            2'b00: ext_data = {24'b0, busRData[7:0]};
                            2'b01: ext_data = {24'b0, busRData[15:8]};
                            2'b10: ext_data = {24'b0, busRData[23:16]};
                            2'b11: ext_data = {24'b0, busRData[31:24]};
                        endcase
                    end
                    3'b101: begin
                        case (half_remain)
                            1'b0: ext_data = {16'b0, busRData[15:0]};
                            1'b1: ext_data = {16'b0, busRData[31:16]};
                        endcase
                    end

                endcase
            end
        endcase
    end
endmodule






module store_bit_concat (
    input  logic [31:0] instrCode,
    input  logic [31:0] RFData2,
    input  logic [31:0] busRData,
    input  logic [31:0] addr,
    output logic [31:0] concat_data
);

    wire [6:0] opcode = instrCode[6:0];
    wire [2:0] func3 = instrCode[14:12];
    wire [1:0] byte_remain = addr[1:0];
    wire half_remain = addr[1];

    always_comb begin
        concat_data = 32'bx;
        case (opcode)
            `OP_TYPE_S: begin
                case (instrCode[14:12])
                    3'b000:
                    case (byte_remain)
                        2'b00: concat_data = {busRData[31:8], RFData2[7:0]};
                        2'b01:
                        concat_data = {
                            busRData[31:16], RFData2[7:0], busRData[7:0]
                        };
                        2'b10:
                        concat_data = {
                            busRData[31:24], RFData2[7:0], busRData[15:0]
                        };
                        2'b11: concat_data = {RFData2[7:0], busRData[23:0]};
                    endcase
                    3'b001:
                    case (half_remain)
                        1'b0: concat_data = {busRData[31:16], RFData2[15:0]};
                        1'b1: concat_data = {RFData2[15:0], busRData[15:0]};
                    endcase
                    3'b010: concat_data = RFData2[31:0];
                endcase
            end
        endcase
    end
endmodule
