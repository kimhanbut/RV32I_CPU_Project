`timescale 1ns / 1ps

module ROM (
    input  logic [31:0] addr,
    output logic [31:0] data
);






  initial begin//////////////////////////// this code for simulation/////////////////////////////////////////////
        $readmemh("code.mem", rom);
        //rom[x]=32'b fucn7 _ rs2 _ rs1 _f3 _ rd  _ op // R-Type
        // rom[0] = 32'b0000000_00001_00010_000_00100_0110011;//add x4, x2, x1
        // rom[1] = 32'b0100000_00001_00011_000_00101_0110011;//sub x5, x3, x1
        // rom[2] = 32'b0000000_00101_10101_001_00110_0110011;//logical left shift x6, x21, x5
        // rom[3] = 32'b0000000_00101_10101_101_00111_0110011;//logical right shift x7, x21, x5

        // rom[4] = 32'b0100000_00001_11111_101_01000_0110011;//arithmetic right shift x8, x31, x1
        // rom[5] = 32'b0100000_00101_10101_101_01001_0110011;//arithmetic right shift x9, x21, x5

        // rom[6] = 32'b0000000_00000_11111_010_01010_0110011;//set less than signed x10, x31, x0
        // rom[7] = 32'b0000000_11111_00000_010_01011_0110011;//set less than signed x11, x0, x31

        // rom[8] = 32'b0000000_00000_11111_011_01100_0110011;//set less than unsigned x12, x31, x0
        // rom[9] = 32'b0000000_11111_00000_011_01101_0110011;//set less than unsigned x13, x0, x31
  end
  assign data = rom[addr[31:2]];


  
    /*/////////////////////////////////////// this code for Design Compiler Synthesis////////////////////////////////////////////
    logic [31:0] word_addr;
    assign word_addr = addr[31:2];
    
    always_comb begin 
        case (word_addr)
            // =====================
            // S-Type: store byte / half
            // =====================
            0:  data = 32'b0000000_11111_00000_000_01111_0100011; // sb x31, 15(x0)
            1:  data = 32'b0000000_11111_00000_000_01110_0100011; // sb x31, 14(x0)
            2:  data = 32'b0000000_11111_00000_000_01101_0100011; // sb x31, 13(x0)
            3:  data = 32'b0000000_11111_00000_001_10110_0100011; // sh x31, 22(x0)
            4:  data = 32'b0000000_11111_00000_001_10100_0100011; // sh x31, 20(x0)

            // =====================
            // L-Type: load byte / half
            // =====================
            5:  data = 32'b0000000_10110_00000_001_01101_0000011; // lh x13, 22(x0)
            6:  data = 32'b0000000_01001_00000_000_01110_0000011; // lb x14, 9(x0)
            7:  data = 32'b0000000_01000_00000_000_01111_0000011; // lb x15, 8(x0)
            8:  data = 32'b0000000_01000_00000_100_10000_0000011; // lbu x16, 8(x0)

            // =====================
            // I-Type
            // =====================
            9:  data = 32'b000000000001_00001_000_01001_0010011; // addi x9, x1, 1
            10: data = 32'b111111111111_00010_000_01010_0010011; // addi x10, x2, -1
            11: data = 32'b000000100000_00011_000_01011_0010011; // addi x11, x3, 32
            12: data = 32'b000000010000_00100_010_01100_0010011; // slti x12, x4, 16
            13: data = 32'b111111111100_00101_010_01101_0010011; // slti x13, x5, -4
            14: data = 32'b000000000001_00110_011_01110_0010011; // sltiu x14, x6, 1
            15: data = 32'b111111111111_00111_011_01111_0010011; // sltiu x15, x7, -1
            16: data = 32'b000000001010_01000_100_10000_0010011; // xori x16, x8, 10
            17: data = 32'b111111110000_01001_100_10001_0010011; // xori x17, x9, -16
            18: data = 32'b000000000111_01010_110_10010_0010011; // ori x18, x10, 7
            19: data = 32'b111111111000_01011_110_10011_0010011; // ori x19, x11, -8
            20: data = 32'b000000001111_01100_111_10100_0010011; // andi x20, x12, 15
            21: data = 32'b111111111111_01101_111_10101_0010011; // andi x21, x13, -1
            22: data = 32'b0000000_00101_01110_001_10110_0010011; // slli x22, x14, 5
            23: data = 32'b0000000_11111_01111_001_10111_0010011; // slli x23, x15, 31
            24: data = 32'b0000000_00101_10000_101_11000_0010011; // srli x24, x16, 5
            25: data = 32'b0100000_00101_10001_101_11001_0010011; // srai x25, x17, 5

            // =====================
            // B-Type: branch (imm = 실제 바이트 이동)
            // =====================

            26: data =32'b0000000_00010_00001_000_01000_1100011;
            27: data =32'b0000000_00011_00001_001_01000_1100011;
            28: data =32'b0000000_00000_00000_000_00000_0000000; 
            29: data =32'b0000000_00100_00001_100_01000_1100011; 
            30: data =32'b0000000_00000_00000_000_01000_0000000; 
            31: data =32'b0000000_00001_00000_101_01000_1100011;
            32: data =32'b0000000_00001_00000_110_01000_1100011; 
            33: data =32'b0000000_00000_00000_000_00000_0000000; 
            34: data =32'b0000000_00000_00001_111_01000_1100011;
            35: data =32'b0000000_00000_00000_000_00000_0000000;

            // =====================
            // LU-Type: LUI
            // =====================
            36: data = 32'b00000000000100100000_00001_0110111;  // LUI x1,0x12000
            37: data = 32'b00000000001101000000_00011_0110111;  // LUI x3,0x34000

            // =====================
            // AU-Type: AUIPC
            // =====================
            38: data = 32'b00000000000100100000_00010_0010111;  // AUIPC x2,0x12000
            39: data = 32'b00000000001101000000_00100_0010111;  // AUIPC x4,0x34000

            // =====================
            // J-Type: JAL (imm = 실제 바이트 이동)
            // =====================
            40: data = {1'b0, 10'd8,9'b0, 5'd5, 7'b1101111}; // JAL x5, +16
            41: data = 32'h00000013; // NOP
            42: data = 32'h00000013; // NOP
            43: data = 32'h00000013; // NOP
            44: data = 32'b00000000101010000000000000010011; // x6 = 42 (JAL target)

            // =====================
            // JALR-Type: JALR (imm = 실제 바이트 이동)
            // =====================
            45: data = 32'b000000001000_00000_000_00111_0010011;  // x7 = 8
            46: data = {12'd200, 5'd7, 3'b000, 5'd8, 7'b1100111};   // JALR x8, x7, 200
            47: data = 32'h00000013; // NOP
            48: data = 32'h00000013; // NOP
            49: data = 32'h00000013; // NOP
            50: data = 32'h00000013; // NOP
            51: data = 32'h00000013; // NOP
            52: data = 32'b0000000110111_00000_000_01001_0010011; // x9 = 55 (JALR target)

            // =====================
            // default: NOP
            // =====================
            default: data = 32'h00000013;  // NOP
        endcase
    end*/
  
endmodule
